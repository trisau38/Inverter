* SPICE3 file created from inverter.ext - technology: scmos

.option scale=1u

M1000 VDD in VDD Gnd nfet w=8 l=2
+  ad=112 pd=72 as=0 ps=0
M1001 VDD in VDD VDD pfet w=24 l=2
+  ad=304 pd=136 as=0 ps=0
C0 VDD Gnd 16.26fF
C1 in Gnd 4.36fF
